`ifndef __CONSTANTS_H__
`define __CONSTANTS_H__

`define SETS 1024
`define TAGS 3
`define WORD_LENGTH 32
`define VALID 1'b1

`define WORD_OFFSET 2
`define ADDR_WORD_OFS_START 1
`define ADDR_WORD_OFS_END 0

`define CACHE_ADDR_LENGTH 10
`define IDX_START 11
`define IDX_END 2

`define CACHE_VALID_BIT 131
`define BLK_TAG_START 130
`define BLK_TAG_END 128

`define TAG_START 14
`define TAG_END 12

`endif